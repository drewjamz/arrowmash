library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Start_Screen_Rom is
    Port (
        addr    : in  STD_LOGIC_VECTOR(13 downto 0); -- 14-bit address input
        data_out: out STD_LOGIC_VECTOR(2 downto 0)  -- 3-bit data output
    );
end Start_Screen_Rom;

architecture Behavioral of Start_Screen_Rom is
begin

    process(addr)
    begin
        case addr is
            when "00000000000000" => data_out <= "000";
            when "00000000000001" => data_out <= "000";
            when "00000000000010" => data_out <= "000";
            when "00000000000011" => data_out <= "000";
            when "00000000000100" => data_out <= "000";
            when "00000000000101" => data_out <= "000";
            when "00000000000110" => data_out <= "000";
            when "00000000000111" => data_out <= "000";
            when "00000000001000" => data_out <= "000";
            when "00000000001001" => data_out <= "000";
            when "00000000001010" => data_out <= "000";
            when "00000000001011" => data_out <= "000";
            when "00000000001100" => data_out <= "000";
            when "00000000001101" => data_out <= "000";
            when "00000000001110" => data_out <= "000";
            when "00000000001111" => data_out <= "000";
            when "00000000010000" => data_out <= "000";
            when "00000000010001" => data_out <= "000";
            when "00000000010010" => data_out <= "000";
            when "00000000010011" => data_out <= "000";
            when "00000000010100" => data_out <= "000";
            when "00000000010101" => data_out <= "000";
            when "00000000010110" => data_out <= "000";
            when "00000000010111" => data_out <= "000";
            when "00000000011000" => data_out <= "000";
            when "00000000011001" => data_out <= "000";
            when "00000000011010" => data_out <= "000";
            when "00000000011011" => data_out <= "000";
            when "00000000011100" => data_out <= "000";
            when "00000000011101" => data_out <= "000";
            when "00000000011110" => data_out <= "000";
            when "00000000011111" => data_out <= "000";
            when "00000000100000" => data_out <= "000";
            when "00000000100001" => data_out <= "000";
            when "00000000100010" => data_out <= "000";
            when "00000000100011" => data_out <= "000";
            when "00000000100100" => data_out <= "000";
            when "00000000100101" => data_out <= "000";
            when "00000000100110" => data_out <= "000";
            when "00000000100111" => data_out <= "000";
            when "00000000101000" => data_out <= "000";
            when "00000000101001" => data_out <= "000";
            when "00000000101010" => data_out <= "000";
            when "00000000101011" => data_out <= "000";
            when "00000000101100" => data_out <= "000";
            when "00000000101101" => data_out <= "000";
            when "00000000101110" => data_out <= "000";
            when "00000000101111" => data_out <= "000";
            when "00000000110000" => data_out <= "000";
            when "00000000110001" => data_out <= "000";
            when "00000000110010" => data_out <= "000";
            when "00000000110011" => data_out <= "000";
            when "00000000110100" => data_out <= "000";
            when "00000000110101" => data_out <= "000";
            when "00000000110110" => data_out <= "000";
            when "00000000110111" => data_out <= "000";
            when "00000000111000" => data_out <= "000";
            when "00000000111001" => data_out <= "000";
            when "00000000111010" => data_out <= "000";
            when "00000000111011" => data_out <= "000";
            when "00000000111100" => data_out <= "000";
            when "00000000111101" => data_out <= "000";
            when "00000000111110" => data_out <= "000";
            when "00000000111111" => data_out <= "000";
            when "00000001000000" => data_out <= "000";
            when "00000001000001" => data_out <= "000";
            when "00000001000010" => data_out <= "000";
            when "00000001000011" => data_out <= "000";
            when "00000001000100" => data_out <= "000";
            when "00000001000101" => data_out <= "000";
            when "00000001000110" => data_out <= "000";
            when "00000001000111" => data_out <= "000";
            when "00000001001000" => data_out <= "000";
            when "00000001001001" => data_out <= "000";
            when "00000001001010" => data_out <= "000";
            when "00000001001011" => data_out <= "000";
            when "00000001001100" => data_out <= "000";
            when "00000001001101" => data_out <= "000";
            when "00000001001110" => data_out <= "000";
            when "00000001001111" => data_out <= "000";
            when "00000001010000" => data_out <= "000";
            when "00000001010001" => data_out <= "000";
            when "00000001010010" => data_out <= "000";
            when "00000001010011" => data_out <= "000";
            when "00000001010100" => data_out <= "000";
            when "00000001010101" => data_out <= "000";
            when "00000001010110" => data_out <= "000";
            when "00000001010111" => data_out <= "000";
            when "00000001011000" => data_out <= "000";
            when "00000001011001" => data_out <= "000";
            when "00000001011010" => data_out <= "000";
            when "00000001011011" => data_out <= "000";
            when "00000001011100" => data_out <= "000";
            when "00000001011101" => data_out <= "000";
            when "00000001011110" => data_out <= "000";
            when "00000001011111" => data_out <= "000";
            when "00000001100000" => data_out <= "000";
            when "00000001100001" => data_out <= "000";
            when "00000001100010" => data_out <= "000";
            when "00000001100011" => data_out <= "000";
            when "00000001100100" => data_out <= "000";
            when "00000001100101" => data_out <= "000";
            when "00000001100110" => data_out <= "000";
            when "00000001100111" => data_out <= "000";
            when "00000001101000" => data_out <= "000";
            when "00000001101001" => data_out <= "000";
            when "00000001101010" => data_out <= "000";
            when "00000001101011" => data_out <= "000";
            when "00000001101100" => data_out <= "000";
            when "00000001101101" => data_out <= "000";
            when "00000001101110" => data_out <= "000";
            when "00000001101111" => data_out <= "000";
            when "00000001110000" => data_out <= "000";
            when "00000001110001" => data_out <= "000";
            when "00000001110010" => data_out <= "000";
            when "00000001110011" => data_out <= "000";
            when "00000001110100" => data_out <= "000";
            when "00000001110101" => data_out <= "000";
            when "00000001110110" => data_out <= "000";
            when "00000001110111" => data_out <= "000";
            when "00000001111000" => data_out <= "000";
            when "00000001111001" => data_out <= "000";
            when "00000001111010" => data_out <= "000";
            when "00000001111011" => data_out <= "000";
            when "00000001111100" => data_out <= "000";
            when "00000001111101" => data_out <= "000";
            when "00000001111110" => data_out <= "000";
            when "00000001111111" => data_out <= "000";
            when "00000010000000" => data_out <= "000";
            when "00000010000001" => data_out <= "000";
            when "00000010000010" => data_out <= "000";
            when "00000010000011" => data_out <= "000";
            when "00000010000100" => data_out <= "000";
            when "00000010000101" => data_out <= "000";
            when "00000010000110" => data_out <= "000";
            when "00000010000111" => data_out <= "000";
            when "00000010001000" => data_out <= "000";
            when "00000010001001" => data_out <= "000";
            when "00000010001010" => data_out <= "000";
            when "00000010001011" => data_out <= "000";
            when "00000010001100" => data_out <= "000";
            when "00000010001101" => data_out <= "000";
            when "00000010001110" => data_out <= "000";
            when "00000010001111" => data_out <= "000";
            when "00000010010000" => data_out <= "000";
            when "00000010010001" => data_out <= "000";
            when "00000010010010" => data_out <= "000";
            when "00000010010011" => data_out <= "000";
            when "00000010010100" => data_out <= "000";
            when "00000010010101" => data_out <= "000";
            when "00000010010110" => data_out <= "000";
            when "00000010010111" => data_out <= "000";
            when "00000010011000" => data_out <= "000";
            when "00000010011001" => data_out <= "000";
            when "00000010011010" => data_out <= "000";
            when "00000010011011" => data_out <= "000";
            when "00000010011100" => data_out <= "000";
            when "00000010011101" => data_out <= "000";
            when "00000010011110" => data_out <= "000";
            when "00000010011111" => data_out <= "000";
            when "00000010100000" => data_out <= "000";
            when "00000010100001" => data_out <= "000";
            when "00000010100010" => data_out <= "000";
            when "00000010100011" => data_out <= "000";
            when "00000010100100" => data_out <= "000";
            when "00000010100101" => data_out <= "000";
            when "00000010100110" => data_out <= "000";
            when "00000010100111" => data_out <= "000";
            when "00000010101000" => data_out <= "000";
            when "00000010101001" => data_out <= "000";
            when "00000010101010" => data_out <= "000";
            when "00000010101011" => data_out <= "000";
            when "00000010101100" => data_out <= "000";
            when "00000010101101" => data_out <= "000";
            when "00000010101110" => data_out <= "000";
            when "00000010101111" => data_out <= "000";
            when "00000010110000" => data_out <= "000";
            when "00000010110001" => data_out <= "000";
            when "00000010110010" => data_out <= "000";
            when "00000010110011" => data_out <= "000";
            when "00000010110100" => data_out <= "000";
            when "00000010110101" => data_out <= "000";
            when "00000010110110" => data_out <= "000";
            when "00000010110111" => data_out <= "000";
            when "00000010111000" => data_out <= "000";
            when "00000010111001" => data_out <= "000";
            when "00000010111010" => data_out <= "000";
            when "00000010111011" => data_out <= "000";
            when "00000010111100" => data_out <= "000";
            when "00000010111101" => data_out <= "000";
            when "00000010111110" => data_out <= "000";
            when "00000010111111" => data_out <= "000";
            when "00000011000000" => data_out <= "000";
            when "00000011000001" => data_out <= "000";
            when "00000011000010" => data_out <= "000";
            when "00000011000011" => data_out <= "000";
            when "00000011000100" => data_out <= "000";
            when "00000011000101" => data_out <= "000";
            when "00000011000110" => data_out <= "000";
            when "00000011000111" => data_out <= "000";
            when "00000011001000" => data_out <= "000";
            when "00000011001001" => data_out <= "000";
            when "00000011001010" => data_out <= "000";
            when "00000011001011" => data_out <= "000";
            when "00000011001100" => data_out <= "000";
            when "00000011001101" => data_out <= "000";
            when "00000011001110" => data_out <= "000";
            when "00000011001111" => data_out <= "000";
            when "00000011010000" => data_out <= "000";
            when "00000011010001" => data_out <= "000";
            when "00000011010010" => data_out <= "000";
            when "00000011010011" => data_out <= "000";
            when "00000011010100" => data_out <= "000";
            when "00000011010101" => data_out <= "000";
            when "00000011010110" => data_out <= "000";
            when "00000011010111" => data_out <= "000";
            when "00000011011000" => data_out <= "000";
            when "00000011011001" => data_out <= "000";
            when "00000011011010" => data_out <= "000";
            when "00000011011011" => data_out <= "000";
            when "00000011011100" => data_out <= "000";
            when "00000011011101" => data_out <= "000";
            when "00000011011110" => data_out <= "000";
            when "00000011011111" => data_out <= "000";
            when "00000011100000" => data_out <= "000";
            when "00000011100001" => data_out <= "000";
            when "00000011100010" => data_out <= "000";
            when "00000011100011" => data_out <= "000";
            when "00000011100100" => data_out <= "000";
            when "00000011100101" => data_out <= "000";
            when "00000011100110" => data_out <= "000";
            when "00000011100111" => data_out <= "000";
            when "00000011101000" => data_out <= "000";
            when "00000011101001" => data_out <= "000";
            when "00000011101010" => data_out <= "000";
            when "00000011101011" => data_out <= "000";
            when "00000011101100" => data_out <= "000";
            when "00000011101101" => data_out <= "000";
            when "00000011101110" => data_out <= "000";
            when "00000011101111" => data_out <= "000";
            when "00000011110000" => data_out <= "000";
            when "00000011110001" => data_out <= "000";
            when "00000011110010" => data_out <= "000";
            when "00000011110011" => data_out <= "000";
            when "00000011110100" => data_out <= "000";
            when "00000011110101" => data_out <= "000";
            when "00000011110110" => data_out <= "000";
            when "00000011110111" => data_out <= "000";
            when "00000011111000" => data_out <= "000";
            when "00000011111001" => data_out <= "000";
            when "00000011111010" => data_out <= "000";
            when "00000011111011" => data_out <= "000";
            when "00000011111100" => data_out <= "000";
            when "00000011111101" => data_out <= "000";
            when "00000011111110" => data_out <= "000";
            when "00000011111111" => data_out <= "000";
            when "00000100000000" => data_out <= "000";
            when "00000100000001" => data_out <= "000";
            when "00000100000010" => data_out <= "000";
            when "00000100000011" => data_out <= "000";
            when "00000100000100" => data_out <= "000";
            when "00000100000101" => data_out <= "000";
            when "00000100000110" => data_out <= "000";
            when "00000100000111" => data_out <= "000";
            when "00000100001000" => data_out <= "000";
            when "00000100001001" => data_out <= "000";
            when "00000100001010" => data_out <= "000";
            when "00000100001011" => data_out <= "000";
            when "00000100001100" => data_out <= "000";
            when "00000100001101" => data_out <= "000";
            when "00000100001110" => data_out <= "000";
            when "00000100001111" => data_out <= "000";
            when "00000100010000" => data_out <= "000";
            when "00000100010001" => data_out <= "000";
            when "00000100010010" => data_out <= "000";
            when "00000100010011" => data_out <= "000";
            when "00000100010100" => data_out <= "000";
            when "00000100010101" => data_out <= "000";
            when "00000100010110" => data_out <= "000";
            when "00000100010111" => data_out <= "000";
            when "00000100011000" => data_out <= "000";
            when "00000100011001" => data_out <= "000";
            when "00000100011010" => data_out <= "000";
            when "00000100011011" => data_out <= "000";
            when "00000100011100" => data_out <= "000";
            when "00000100011101" => data_out <= "000";
            when "00000100011110" => data_out <= "000";
            when "00000100011111" => data_out <= "000";
            when "00000100100000" => data_out <= "000";
            when "00000100100001" => data_out <= "000";
            when "00000100100010" => data_out <= "000";
            when "00000100100011" => data_out <= "000";
            when "00000100100100" => data_out <= "000";
            when "00000100100101" => data_out <= "000";
            when "00000100100110" => data_out <= "000";
            when "00000100100111" => data_out <= "000";
            when "00000100101000" => data_out <= "000";
            when "00000100101001" => data_out <= "000";
            when "00000100101010" => data_out <= "000";
            when "00000100101011" => data_out <= "000";
            when "00000100101100" => data_out <= "000";
            when "00000100101101" => data_out <= "000";
            when "00000100101110" => data_out <= "000";
            when "00000100101111" => data_out <= "000";
            when "00000100110000" => data_out <= "000";
            when "00000100110001" => data_out <= "000";
            when "00000100110010" => data_out <= "000";
            when "00000100110011" => data_out <= "000";
            when "00000100110100" => data_out <= "000";
            when "00000100110101" => data_out <= "000";
            when "00000100110110" => data_out <= "000";
            when "00000100110111" => data_out <= "000";
            when "00000100111000" => data_out <= "000";
            when "00000100111001" => data_out <= "000";
            when "00000100111010" => data_out <= "000";
            when "00000100111011" => data_out <= "000";
            when "00000100111100" => data_out <= "000";
            when "00000100111101" => data_out <= "000";
            when "00000100111110" => data_out <= "000";
            when "00000100111111" => data_out <= "000";
            when "00000101000000" => data_out <= "000";
            when "00000101000001" => data_out <= "000";
            when "00000101000010" => data_out <= "000";
            when "00000101000011" => data_out <= "000";
            when "00000101000100" => data_out <= "000";
            when "00000101000101" => data_out <= "000";
            when "00000101000110" => data_out <= "000";
            when "00000101000111" => data_out <= "000";
            when "00000101001000" => data_out <= "000";
            when "00000101001001" => data_out <= "000";
            when "00000101001010" => data_out <= "000";
            when "00000101001011" => data_out <= "000";
            when "00000101001100" => data_out <= "000";
            when "00000101001101" => data_out <= "000";
            when "00000101001110" => data_out <= "000";
            when "00000101001111" => data_out <= "000";
            when "00000101010000" => data_out <= "000";
            when "00000101010001" => data_out <= "000";
            when "00000101010010" => data_out <= "000";
            when "00000101010011" => data_out <= "000";
            when "00000101010100" => data_out <= "000";
            when "00000101010101" => data_out <= "000";
            when "00000101010110" => data_out <= "000";
            when "00000101010111" => data_out <= "000";
            when "00000101011000" => data_out <= "000";
            when "00000101011001" => data_out <= "000";
            when "00000101011010" => data_out <= "000";
            when "00000101011011" => data_out <= "000";
            when "00000101011100" => data_out <= "000";
            when "00000101011101" => data_out <= "000";
            when "00000101011110" => data_out <= "000";
            when "00000101011111" => data_out <= "000";
            when "00000101100000" => data_out <= "000";
            when "00000101100001" => data_out <= "000";
            when "00000101100010" => data_out <= "000";
            when "00000101100011" => data_out <= "000";
            when "00000101100100" => data_out <= "000";
            when "00000101100101" => data_out <= "000";
            when "00000101100110" => data_out <= "000";
            when "00000101100111" => data_out <= "000";
            when "00000101101000" => data_out <= "000";
            when "00000101101001" => data_out <= "000";
            when "00000101101010" => data_out <= "000";
            when "00000101101011" => data_out <= "000";
            when "00000101101100" => data_out <= "000";
            when "00000101101101" => data_out <= "000";
            when "00000101101110" => data_out <= "000";
            when "00000101101111" => data_out <= "000";
            when "00000101110000" => data_out <= "000";
            when "00000101110001" => data_out <= "000";
            when "00000101110010" => data_out <= "000";
            when "00000101110011" => data_out <= "000";
            when "00000101110100" => data_out <= "000";
            when "00000101110101" => data_out <= "000";
            when "00000101110110" => data_out <= "000";
            when "00000101110111" => data_out <= "000";
            when "00000101111000" => data_out <= "000";
            when "00000101111001" => data_out <= "000";
            when "00000101111010" => data_out <= "000";
            when "00000101111011" => data_out <= "000";
            when "00000101111100" => data_out <= "000";
            when "00000101111101" => data_out <= "000";
            when "00000101111110" => data_out <= "000";
            when "00000101111111" => data_out <= "000";
            when "00000110000000" => data_out <= "000";
            when "00000110000001" => data_out <= "000";
            when "00000110000010" => data_out <= "000";
            when "00000110000011" => data_out <= "000";
            when "00000110000100" => data_out <= "000";
            when "00000110000101" => data_out <= "000";
            when "00000110000110" => data_out <= "000";
            when "00000110000111" => data_out <= "000";
            when "00000110001000" => data_out <= "000";
            when "00000110001001" => data_out <= "000";
            when "00000110001010" => data_out <= "000";
            when "00000110001011" => data_out <= "000";
            when "00000110001100" => data_out <= "000";
            when "00000110001101" => data_out <= "000";
            when "00000110001110" => data_out <= "000";
            when "00000110001111" => data_out <= "000";
            when "00000110010000" => data_out <= "000";
            when "00000110010001" => data_out <= "000";
            when "00000110010010" => data_out <= "000";
            when "00000110010011" => data_out <= "000";
            when "00000110010100" => data_out <= "000";
            when "00000110010101" => data_out <= "000";
            when "00000110010110" => data_out <= "000";
            when "00000110010111" => data_out <= "000";
            when "00000110011000" => data_out <= "000";
            when "00000110011001" => data_out <= "000";
            when "00000110011010" => data_out <= "000";
            when "00000110011011" => data_out <= "000";
            when "00000110011100" => data_out <= "000";
            when "00000110011101" => data_out <= "000";
            when "00000110011110" => data_out <= "000";
            when "00000110011111" => data_out <= "000";
            when "00000110100000" => data_out <= "000";
            when "00000110100001" => data_out <= "000";
            when "00000110100010" => data_out <= "000";
            when "00000110100011" => data_out <= "000";
            when "00000110100100" => data_out <= "000";
            when "00000110100101" => data_out <= "000";
            when "00000110100110" => data_out <= "000";
            when "00000110100111" => data_out <= "000";
            when "00000110101000" => data_out <= "000";
            when "00000110101001" => data_out <= "000";
            when "00000110101010" => data_out <= "000";
            when "00000110101011" => data_out <= "000";
            when "00000110101100" => data_out <= "000";
            when "00000110101101" => data_out <= "000";
            when "00000110101110" => data_out <= "000";
            when "00000110101111" => data_out <= "000";
            when "00000110110000" => data_out <= "000";
            when "00000110110001" => data_out <= "000";
            when "00000110110010" => data_out <= "000";
            when "00000110110011" => data_out <= "000";
            when "00000110110100" => data_out <= "000";
            when "00000110110101" => data_out <= "000";
            when "00000110110110" => data_out <= "000";
            when "00000110110111" => data_out <= "000";
            when "00000110111000" => data_out <= "000";
            when "00000110111001" => data_out <= "000";
            when "00000110111010" => data_out <= "000";
            when "00000110111011" => data_out <= "000";
            when "00000110111100" => data_out <= "000";
            when "00000110111101" => data_out <= "000";
            when "00000110111110" => data_out <= "000";
            when "00000110111111" => data_out <= "000";
            when "00000111000000" => data_out <= "000";
            when "00000111000001" => data_out <= "000";
            when "00000111000010" => data_out <= "000";
            when "00000111000011" => data_out <= "000";
            when "00000111000100" => data_out <= "000";
            when "00000111000101" => data_out <= "000";
            when "00000111000110" => data_out <= "000";
            when "00000111000111" => data_out <= "000";
            when "00000111001000" => data_out <= "000";
            when "00000111001001" => data_out <= "000";
            when "00000111001010" => data_out <= "000";
            when "00000111001011" => data_out <= "000";
            when "00000111001100" => data_out <= "000";
            when "00000111001101" => data_out <= "000";
            when "00000111001110" => data_out <= "000";
            when "00000111001111" => data_out <= "000";
            when "00000111010000" => data_out <= "000";
            when "00000111010001" => data_out <= "000";
            when "00000111010010" => data_out <= "000";
            when "00000111010011" => data_out <= "000";
            when "00000111010100" => data_out <= "000";
            when "00000111010101" => data_out <= "000";
            when "00000111010110" => data_out <= "000";
            when "00000111010111" => data_out <= "000";
            when "00000111011000" => data_out <= "000";
            when "00000111011001" => data_out <= "000";
            when "00000111011010" => data_out <= "000";
            when "00000111011011" => data_out <= "000";
            when "00000111011100" => data_out <= "000";
            when "00000111011101" => data_out <= "000";
            when "00000111011110" => data_out <= "000";
            when "00000111011111" => data_out <= "000";
            when "00000111100000" => data_out <= "000";
            when "00000111100001" => data_out <= "000";
            when "00000111100010" => data_out <= "000";
            when "00000111100011" => data_out <= "000";
            when "00000111100100" => data_out <= "000";
            when "00000111100101" => data_out <= "000";
            when "00000111100110" => data_out <= "000";
            when "00000111100111" => data_out <= "000";
            when "00000111101000" => data_out <= "000";
            when "00000111101001" => data_out <= "000";
            when "00000111101010" => data_out <= "000";
            when "00000111101011" => data_out <= "000";
            when "00000111101100" => data_out <= "000";
            when "00000111101101" => data_out <= "000";
            when "00000111101110" => data_out <= "000";
            when "00000111101111" => data_out <= "000";
            when "00000111110000" => data_out <= "000";
            when "00000111110001" => data_out <= "000";
            when "00000111110010" => data_out <= "000";
            when "00000111110011" => data_out <= "000";
            when "00000111110100" => data_out <= "000";
            when "00000111110101" => data_out <= "000";
            when "00000111110110" => data_out <= "000";
            when "00000111110111" => data_out <= "000";
            when "00000111111000" => data_out <= "000";
            when "00000111111001" => data_out <= "000";
            when "00000111111010" => data_out <= "000";
            when "00000111111011" => data_out <= "000";
            when "00000111111100" => data_out <= "000";
            when "00000111111101" => data_out <= "000";
            when "00000111111110" => data_out <= "000";
            when "00000111111111" => data_out <= "000";
            when "00001000000000" => data_out <= "000";
            when "00001000000001" => data_out <= "000";
            when "00001000000010" => data_out <= "000";
            when "00001000000011" => data_out <= "000";
            when "00001000000100" => data_out <= "000";
            when "00001000000101" => data_out <= "000";
            when "00001000000110" => data_out <= "000";
            when "00001000000111" => data_out <= "000";
            when "00001000001000" => data_out <= "000";
            when "00001000001001" => data_out <= "000";
            when "00001000001010" => data_out <= "000";
            when "00001000001011" => data_out <= "000";
            when "00001000001100" => data_out <= "000";
            when "00001000001101" => data_out <= "000";
            when "00001000001110" => data_out <= "000";
            when "00001000001111" => data_out <= "000";
            when "00001000010000" => data_out <= "000";
            when "00001000010001" => data_out <= "000";
            when "00001000010010" => data_out <= "000";
            when "00001000010011" => data_out <= "000";
            when "00001000010100" => data_out <= "000";
            when "00001000010101" => data_out <= "000";
            when "00001000010110" => data_out <= "000";
            when "00001000010111" => data_out <= "000";
            when "00001000011000" => data_out <= "000";
            when "00001000011001" => data_out <= "000";
            when "00001000011010" => data_out <= "000";
            when "00001000011011" => data_out <= "000";
            when "00001000011100" => data_out <= "000";
            when "00001000011101" => data_out <= "000";
            when "00001000011110" => data_out <= "000";
            when "00001000011111" => data_out <= "000";
            when "00001000100000" => data_out <= "111";
            when "00001000100001" => data_out <= "111";
            when "00001000100010" => data_out <= "111";
            when "00001000100011" => data_out <= "111";
            when "00001000100100" => data_out <= "111";
            when "00001000100101" => data_out <= "111";
            when "00001000100110" => data_out <= "111";
            when "00001000100111" => data_out <= "111";
            when "00001000101000" => data_out <= "111";
            when "00001000101001" => data_out <= "111";
            when "00001000101010" => data_out <= "111";
            when "00001000101011" => data_out <= "111";
            when "00001000101100" => data_out <= "111";
            when "00001000101101" => data_out <= "111";
            when "00001000101110" => data_out <= "111";
            when "00001000101111" => data_out <= "111";
            when "00001000110000" => data_out <= "111";
            when "00001000110001" => data_out <= "111";
            when "00001000110010" => data_out <= "111";
            when "00001000110011" => data_out <= "111";
            when "00001000110100" => data_out <= "111";
            when "00001000110101" => data_out <= "111";
            when "00001000110110" => data_out <= "000";
            when "00001000110111" => data_out <= "000";
            when "00001000111000" => data_out <= "000";
            when "00001000111001" => data_out <= "000";
            when "00001000111010" => data_out <= "000";
            when "00001000111011" => data_out <= "000";
            when "00001000111100" => data_out <= "000";
            when "00001000111101" => data_out <= "000";
            when "00001000111110" => data_out <= "000";
            when "00001000111111" => data_out <= "000";
            when "00001001000000" => data_out <= "000";
            when "00001001000001" => data_out <= "000";
            when "00001001000010" => data_out <= "000";
            when "00001001000011" => data_out <= "000";
            when "00001001000100" => data_out <= "000";
            when "00001001000101" => data_out <= "000";
            when "00001001000110" => data_out <= "000";
            when "00001001000111" => data_out <= "000";
            when "00001001001000" => data_out <= "000";
            when "00001001001001" => data_out <= "000";
            when "00001001001010" => data_out <= "000";
            when "00001001001011" => data_out <= "000";
            when "00001001001100" => data_out <= "000";
            when "00001001001101" => data_out <= "000";
            when "00001001001110" => data_out <= "111";
            when "00001001001111" => data_out <= "000";
            when "00001001010000" => data_out <= "111";
            when "00001001010001" => data_out <= "111";
            when "00001001010010" => data_out <= "000";
            when "00001001010011" => data_out <= "000";
            when "00001001010100" => data_out <= "000";
            when "00001001010101" => data_out <= "000";
            when "00001001010110" => data_out <= "000";
            when "00001001010111" => data_out <= "000";
            when "00001001011000" => data_out <= "000";
            when "00001001011001" => data_out <= "000";
            when "00001001011010" => data_out <= "000";
            when "00001001011011" => data_out <= "000";
            when "00001001011100" => data_out <= "000";
            when "00001001011101" => data_out <= "000";
            when "00001001011110" => data_out <= "000";
            when "00001001011111" => data_out <= "000";
            when "00001001100000" => data_out <= "000";
            when "00001001100001" => data_out <= "000";
            when "00001001100010" => data_out <= "000";
            when "00001001100011" => data_out <= "000";
            when "00001001100100" => data_out <= "000";
            when "00001001100101" => data_out <= "000";
            when "00001001100110" => data_out <= "000";
            when "00001001100111" => data_out <= "000";
            when "00001001101000" => data_out <= "000";
            when "00001001101001" => data_out <= "000";
            when "00001001101010" => data_out <= "000";
            when "00001001101011" => data_out <= "000";
            when "00001001101100" => data_out <= "000";
            when "00001001101101" => data_out <= "000";
            when "00001001101110" => data_out <= "000";
            when "00001001101111" => data_out <= "000";
            when "00001001110000" => data_out <= "000";
            when "00001001110001" => data_out <= "000";
            when "00001001110010" => data_out <= "000";
            when "00001001110011" => data_out <= "000";
            when "00001001110100" => data_out <= "000";
            when "00001001110101" => data_out <= "000";
            when "00001001110110" => data_out <= "000";
            when "00001001110111" => data_out <= "000";
            when "00001001111000" => data_out <= "000";
            when "00001001111001" => data_out <= "000";
            when "00001001111010" => data_out <= "000";
            when "00001001111011" => data_out <= "000";
            when "00001001111100" => data_out <= "000";
            when "00001001111101" => data_out <= "000";
            when "00001001111110" => data_out <= "000";
            when "00001001111111" => data_out <= "000";
            when "00001010000000" => data_out <= "000";
            when "00001010000001" => data_out <= "000";
            when "00001010000010" => data_out <= "000";
            when "00001010000011" => data_out <= "000";
            when "00001010000100" => data_out <= "000";
            when "00001010000101" => data_out <= "000";
            when "00001010000110" => data_out <= "000";
            when "00001010000111" => data_out <= "000";
            when "00001010001000" => data_out <= "000";
            when "00001010001001" => data_out <= "000";
            when "00001010001010" => data_out <= "000";
            when "00001010001011" => data_out <= "000";
            when "00001010001100" => data_out <= "000";
            when "00001010001101" => data_out <= "000";
            when "00001010001110" => data_out <= "000";
            when "00001010001111" => data_out <= "000";
            when "00001010010000" => data_out <= "000";
            when "00001010010001" => data_out <= "000";
            when "00001010010010" => data_out <= "000";
            when "00001010010011" => data_out <= "000";
            when "00001010010100" => data_out <= "000";
            when "00001010010101" => data_out <= "000";
            when "00001010010110" => data_out <= "000";
            when "00001010010111" => data_out <= "000";
            when "00001010011000" => data_out <= "000";
            when "00001010011001" => data_out <= "000";
            when "00001010011010" => data_out <= "000";
            when "00001010011011" => data_out <= "000";
            when "00001010011100" => data_out <= "111";
            when "00001010011101" => data_out <= "111";
            when "00001010011110" => data_out <= "111";
            when "00001010011111" => data_out <= "111";
            when "00001010100000" => data_out <= "100";
            when "00001010100001" => data_out <= "100";
            when "00001010100010" => data_out <= "000";
            when "00001010100011" => data_out <= "100";
            when "00001010100100" => data_out <= "100";
            when "00001010100101" => data_out <= "000";
            when "00001010100110" => data_out <= "100";
            when "00001010100111" => data_out <= "100";
            when "00001010101000" => data_out <= "100";
            when "00001010101001" => data_out <= "100";
            when "00001010101010" => data_out <= "100";
            when "00001010101011" => data_out <= "100";
            when "00001010101100" => data_out <= "100";
            when "00001010101101" => data_out <= "100";
            when "00001010101110" => data_out <= "100";
            when "00001010101111" => data_out <= "100";
            when "00001010110000" => data_out <= "100";
            when "00001010110001" => data_out <= "100";
            when "00001010110010" => data_out <= "111";
            when "00001010110011" => data_out <= "111";
            when "00001010110100" => data_out <= "111";
            when "00001010110101" => data_out <= "111";
            when "00001010110110" => data_out <= "000";
            when "00001010110111" => data_out <= "000";
            when "00001010111000" => data_out <= "000";
            when "00001010111001" => data_out <= "000";
            when "00001010111010" => data_out <= "000";
            when "00001010111011" => data_out <= "000";
            when "00001010111100" => data_out <= "000";
            when "00001010111101" => data_out <= "000";
            when "00001010111110" => data_out <= "000";
            when "00001010111111" => data_out <= "000";
            when "00001011000000" => data_out <= "000";
            when "00001011000001" => data_out <= "000";
            when "00001011000010" => data_out <= "000";
            when "00001011000011" => data_out <= "000";
            when "00001011000100" => data_out <= "000";
            when "00001011000101" => data_out <= "000";
            when "00001011000110" => data_out <= "000";
            when "00001011000111" => data_out <= "000";
            when "00001011001000" => data_out <= "000";
            when "00001011001001" => data_out <= "000";
            when "00001011001010" => data_out <= "000";
            when "00001011001011" => data_out <= "000";
            when "00001011001100" => data_out <= "000";
            when "00001011001101" => data_out <= "000";
            when "00001011001110" => data_out <= "000";
            when "00001011001111" => data_out <= "000";
            when "00001011010000" => data_out <= "111";
            when "00001011010001" => data_out <= "111";
            when "00001011010010" => data_out <= "111";
            when "00001011010011" => data_out <= "111";
            when "00001011010100" => data_out <= "111";
            when "00001011010101" => data_out <= "111";
            when "00001011010110" => data_out <= "000";
            when "00001011010111" => data_out <= "000";
            when "00001011011000" => data_out <= "000";
            when "00001011011001" => data_out <= "000";
            when "00001011011010" => data_out <= "000";
            when "00001011011011" => data_out <= "000";
            when "00001011011100" => data_out <= "000";
            when "00001011011101" => data_out <= "000";
            when "00001011011110" => data_out <= "000";
            when "00001011011111" => data_out <= "000";
            when "00001011100000" => data_out <= "000";
            when "00001011100001" => data_out <= "000";
            when "00001011100010" => data_out <= "000";
            when "00001011100011" => data_out <= "000";
            when "00001011100100" => data_out <= "000";
            when "00001011100101" => data_out <= "000";
            when "00001011100110" => data_out <= "000";
            when "00001011100111" => data_out <= "000";
            when "00001011101000" => data_out <= "000";
            when "00001011101001" => data_out <= "000";
            when "00001011101010" => data_out <= "000";
            when "00001011101011" => data_out <= "000";
            when "00001011101100" => data_out <= "000";
            when "00001011101101" => data_out <= "000";
            when "00001011101110" => data_out <= "000";
            when "00001011101111" => data_out <= "000";
            when "00001011110000" => data_out <= "000";
            when "00001011110001" => data_out <= "000";
            when "00001011110010" => data_out <= "000";
            when "00001011110011" => data_out <= "000";
            when "00001011110100" => data_out <= "000";
            when "00001011110101" => data_out <= "000";
            when "00001011110110" => data_out <= "000";
            when "00001011110111" => data_out <= "000";
            when "00001011111000" => data_out <= "000";
            when "00001011111001" => data_out <= "000";
            when "00001011111010" => data_out <= "000";
            when "00001011111011" => data_out <= "000";
            when "00001011111100" => data_out <= "000";
            when "00001011111101" => data_out <= "000";
            when "00001011111110" => data_out <= "000";
            when "00001011111111" => data_out <= "000";
            when "00001100000000" => data_out <= "000";
            when "00001100000001" => data_out <= "000";
            when "00001100000010" => data_out <= "000";
            when "00001100000011" => data_out <= "000";
            when "00001100000100" => data_out <= "000";
            when "00001100000101" => data_out <= "000";
            when "00001100000110" => data_out <= "000";
            when "00001100000111" => data_out <= "000";
            when "00001100001000" => data_out <= "000";
            when "00001100001001" => data_out <= "000";
            when "00001100001010" => data_out <= "000";
            when "00001100001011" => data_out <= "000";
            when "00001100001100" => data_out <= "000";
            when "00001100001101" => data_out <= "000";
            when "00001100001110" => data_out <= "000";
            when "00001100001111" => data_out <= "000";
            when "00001100010000" => data_out <= "000";
            when "00001100010001" => data_out <= "000";
            when "00001100010010" => data_out <= "000";
            when "00001100010011" => data_out <= "000";
            when "00001100010100" => data_out <= "000";
            when "00001100010101" => data_out <= "000";
            when "00001100010110" => data_out <= "000";
            when "00001100010111" => data_out <= "000";
            when "00001100011000" => data_out <= "000";
            when "00001100011001" => data_out <= "000";
            when "00001100011010" => data_out <= "000";
            when "00001100011011" => data_out <= "000";
            when "00001100011100" => data_out <= "111";
            when "00001100011101" => data_out <= "111";
            when "00001100011110" => data_out <= "111";
            when "00001100011111" => data_out <= "111";
            when "00001100100000" => data_out <= "100";
            when "00001100100001" => data_out <= "100";
            when "00001100100010" => data_out <= "000";
            when "00001100100011" => data_out <= "100";
            when "00001100100100" => data_out <= "100";
            when "00001100100101" => data_out <= "000";
            when "00001100100110" => data_out <= "000";
            when "00001100100111" => data_out <= "100";
            when "00001100101000" => data_out <= "100";
            when "00001100101001" => data_out <= "100";
            when "00001100101010" => data_out <= "100";
            when "00001100101011" => data_out <= "100";
            when "00001100101100" => data_out <= "000";
            when "00001100101101" => data_out <= "100";
            when "00001100101110" => data_out <= "100";
            when "00001100101111" => data_out <= "100";
            when "00001100110000" => data_out <= "100";
            when "00001100110001" => data_out <= "100";
            when "00001100110010" => data_out <= "111";
            when "00001100110011" => data_out <= "111";
            when "00001100110100" => data_out <= "111";
            when "00001100110101" => data_out <= "111";
            when "00001100110110" => data_out <= "000";
            when "00001100110111" => data_out <= "000";
            when "00001100111000" => data_out <= "000";
            when "00001100111001" => data_out <= "000";
            when "00001100111010" => data_out <= "000";
            when "00001100111011" => data_out <= "000";
            when "00001100111100" => data_out <= "000";
            when "00001100111101" => data_out <= "000";
            when "00001100111110" => data_out <= "000";
            when "00001100111111" => data_out <= "000";
            when "00001101000000" => data_out <= "000";
            when "00001101000001" => data_out <= "000";
            when "00001101000010" => data_out <= "000";
            when "00001101000011" => data_out <= "000";
            when "00001101000100" => data_out <= "000";
            when "00001101000101" => data_out <= "000";
            when "00001101000110" => data_out <= "000";
            when "00001101000111" => data_out <= "000";
            when "00001101001000" => data_out <= "000";
            when "00001101001001" => data_out <= "000";
            when "00001101001010" => data_out <= "000";
            when "00001101001011" => data_out <= "000";
            when "00001101001100" => data_out <= "000";
            when "00001101001101" => data_out <= "000";
            when "00001101001110" => data_out <= "111";
            when "00001101001111" => data_out <= "000";
            when "00001101010000" => data_out <= "000";
            when "00001101010001" => data_out <= "111";
            when "00001101010010" => data_out <= "000";
            when "00001101010011" => data_out <= "000";
            when "00001101010100" => data_out <= "000";
            when "00001101010101" => data_out <= "111";
            when "00001101010110" => data_out <= "000";
            when "00001101010111" => data_out <= "000";
            when "00001101011000" => data_out <= "000";
            when "00001101011001" => data_out <= "000";
            when "00001101011010" => data_out <= "000";
            when "00001101011011" => data_out <= "000";
            when "00001101011100" => data_out <= "000";
            when "00001101011101" => data_out <= "000";
            when "00001101011110" => data_out <= "000";
            when "00001101011111" => data_out <= "000";
            when "00001101100000" => data_out <= "000";
            when "00001101100001" => data_out <= "000";
            when "00001101100010" => data_out <= "000";
            when "00001101100011" => data_out <= "000";
            when "00001101100100" => data_out <= "000";
            when "00001101100101" => data_out <= "000";
            when "00001101100110" => data_out <= "000";
            when "00001101100111" => data_out <= "000";
            when "00001101101000" => data_out <= "000";
            when "00001101101001" => data_out <= "000";
            when "00001101101010" => data_out <= "000";
            when "00001101101011" => data_out <= "000";
            when "00001101101100" => data_out <= "000";
            when "00001101101101" => data_out <= "000";
            when "00001101101110" => data_out <= "000";
            when "00001101101111" => data_out <= "000";
            when "00001101110000" => data_out <= "000";
            when "00001101110001" => data_out <= "000";
            when "00001101110010" => data_out <= "000";
            when "00001101110011" => data_out <= "000";
            when "00001101110100" => data_out <= "000";
            when "00001101110101" => data_out <= "000";
            when "00001101110110" => data_out <= "000";
            when "00001101110111" => data_out <= "000";
            when "00001101111000" => data_out <= "000";
            when "00001101111001" => data_out <= "000";
            when "00001101111010" => data_out <= "000";
            when "00001101111011" => data_out <= "000";
            when "00001101111100" => data_out <= "000";
            when "00001101111101" => data_out <= "000";
            when "00001101111110" => data_out <= "000";
            when "00001101111111" => data_out <= "000";
            when "00001110000000" => data_out <= "000";
            when "00001110000001" => data_out <= "000";
            when "00001110000010" => data_out <= "000";
            when "00001110000011" => data_out <= "000";
            when "00001110000100" => data_out <= "000";
            when "00001110000101" => data_out <= "000";
            when "00001110000110" => data_out <= "000";
            when "00001110000111" => data_out <= "000";
            when "00001110001000" => data_out <= "000";
            when "00001110001001" => data_out <= "000";
            when "00001110001010" => data_out <= "000";
            when "00001110001011" => data_out <= "000";
            when "00001110001100" => data_out <= "000";
            when "00001110001101" => data_out <= "000";
            when "00001110001110" => data_out <= "000";
            when "00001110001111" => data_out <= "000";
            when "00001110010000" => data_out <= "000";
            when "00001110010001" => data_out <= "000";
            when "00001110010010" => data_out <= "000";
            when "00001110010011" => data_out <= "000";
            when "00001110010100" => data_out <= "000";
            when "00001110010101" => data_out <= "000";
            when "00001110010110" => data_out <= "000";
            when "00001110010111" => data_out <= "000";
            when "00001110011000" => data_out <= "000";
            when "00001110011001" => data_out <= "000";
            when "00001110011010" => data_out <= "000";
            when "00001110011011" => data_out <= "000";
            when "00001110011100" => data_out <= "111";
            when "00001110011101" => data_out <= "111";
            when "00001110011110" => data_out <= "111";
            when "00001110011111" => data_out <= "111";
            when "00001110100000" => data_out <= "100";
            when "00001110100001" => data_out <= "100";
            when "00001110100010" => data_out <= "100";
            when "00001110100011" => data_out <= "100";
            when "00001110100100" => data_out <= "100";
            when "00001110100101" => data_out <= "100";
            when "00001110100110" => data_out <= "100";
            when "00001110100111" => data_out <= "100";
            when "00001110101000" => data_out <= "100";
            when "00001110101001" => data_out <= "100";
            when "00001110101010" => data_out <= "000";
            when "00001110101011" => data_out <= "100";
            when "00001110101100" => data_out <= "100";
            when "00001110101101" => data_out <= "000";
            when "00001110101110" => data_out <= "100";
            when "00001110101111" => data_out <= "100";
            when "00001110110000" => data_out <= "100";
            when "00001110110001" => data_out <= "100";
            when "00001110110010" => data_out <= "111";
            when "00001110110011" => data_out <= "111";
            when "00001110110100" => data_out <= "111";
            when "00001110110101" => data_out <= "111";
            when "00001110110110" => data_out <= "000";
            when "00001110110111" => data_out <= "000";
            when "00001110111000" => data_out <= "000";
            when "00001110111001" => data_out <= "000";
            when "00001110111010" => data_out <= "000";
            when "00001110111011" => data_out <= "000";
            when "00001110111100" => data_out <= "000";
            when "00001110111101" => data_out <= "000";
            when "00001110111110" => data_out <= "000";
            when "00001110111111" => data_out <= "000";
            when "00001111000000" => data_out <= "000";
            when "00001111000001" => data_out <= "000";
            when "00001111000010" => data_out <= "000";
            when "00001111000011" => data_out <= "000";
            when "00001111000100" => data_out <= "000";
            when "00001111000101" => data_out <= "000";
            when "00001111000110" => data_out <= "000";
            when "00001111000111" => data_out <= "000";
            when "00001111001000" => data_out <= "000";
            when "00001111001001" => data_out <= "000";
            when "00001111001010" => data_out <= "000";
            when "00001111001011" => data_out <= "000";
            when "00001111001100" => data_out <= "000";
            when "00001111001101" => data_out <= "000";
            when "00001111001110" => data_out <= "111";
            when "00001111001111" => data_out <= "000";
            when "00001111010000" => data_out <= "000";
            when "00001111010001" => data_out <= "111";
            when "00001111010010" => data_out <= "111";
            when "00001111010011" => data_out <= "111";
            when "00001111010100" => data_out <= "111";
            when "00001111010101" => data_out <= "111";
            when "00001111010110" => data_out <= "000";
            when "00001111010111" => data_out <= "000";
            when "00001111011000" => data_out <= "000";
            when "00001111011001" => data_out <= "000";
            when "00001111011010" => data_out <= "000";
            when "00001111011011" => data_out <= "000";
            when "00001111011100" => data_out <= "000";
            when "00001111011101" => data_out <= "000";
            when "00001111011110" => data_out <= "000";
            when "00001111011111" => data_out <= "000";
            when "00001111100000" => data_out <= "000";
            when "00001111100001" => data_out <= "000";
            when "00001111100010" => data_out <= "000";
            when "00001111100011" => data_out <= "000";
            when "00001111100100" => data_out <= "000";
            when "00001111100101" => data_out <= "000";
            when "00001111100110" => data_out <= "000";
            when "00001111100111" => data_out <= "000";
            when "00001111101000" => data_out <= "000";
            when "00001111101001" => data_out <= "000";
            when "00001111101010" => data_out <= "000";
            when "00001111101011" => data_out <= "000";
            when "00001111101100" => data_out <= "000";
            when "00001111101101" => data_out <= "000";
            when "00001111101110" => data_out <= "000";
            when "00001111101111" => data_out <= "000";
            when "00001111110000" => data_out <= "000";
            when "00001111110001" => data_out <= "000";
            when "00001111110010" => data_out <= "000";
            when "00001111110011" => data_out <= "000";
            when "00001111110100" => data_out <= "000";
            when "00001111110101" => data_out <= "000";
            when "00001111110110" => data_out <= "000";
            when "00001111110111" => data_out <= "000";
            when "00001111111000" => data_out <= "000";
            when "00001111111001" => data_out <= "000";
            when "00001111111010" => data_out <= "000";
            when "00001111111011" => data_out <= "000";
            when "00001111111100" => data_out <= "000";
            when "00001111111101" => data_out <= "000";
            when "00001111111110" => data_out <= "000";
            when "00001111111111" => data_out <= "000";
            when "00010000000000" => data_out <= "000";
            when "00010000000001" => data_out <= "000";
            when "00010000000010" => data_out <= "000";
            when "00010000000011" => data_out <= "000";
            when "00010000000100" => data_out <= "000";
            when "00010000000101" => data_out <= "000";
            when "00010000000110" => data_out <= "000";
            when "00010000000111" => data_out <= "000";
            when "00010000001000" => data_out <= "000";
            when "00010000001001" => data_out <= "000";
            when "00010000001010" => data_out <= "000";
            when "00010000001011" => data_out <= "000";
            when "00010000001100" => data_out <= "000";
            when "00010000001101" => data_out <= "000";
            when "00010000001110" => data_out <= "000";
            when "00010000001111" => data_out <= "000";
            when "00010000010000" => data_out <= "000";
            when "00010000010001" => data_out <= "000";
            when "00010000010010" => data_out <= "000";
            when "00010000010011" => data_out <= "000";
            when "00010000010100" => data_out <= "000";
            when "00010000010101" => data_out <= "000";
            when "00010000010110" => data_out <= "000";
            when "00010000010111" => data_out <= "000";
            when "00010000011000" => data_out <= "000";
            when "00010000011001" => data_out <= "000";
            when "00010000011010" => data_out <= "000";
            when "00010000011011" => data_out <= "000";
            when "00010000011100" => data_out <= "111";
            when "00010000011101" => data_out <= "111";
            when "00010000011110" => data_out <= "111";
            when "00010000011111" => data_out <= "111";
            when "00010000100000" => data_out <= "100";
            when "00010000100001" => data_out <= "100";
            when "00010000100010" => data_out <= "100";
            when "00010000100011" => data_out <= "100";
            when "00010000100100" => data_out <= "000";
            when "00010000100101" => data_out <= "000";
            when "00010000100110" => data_out <= "100";
            when "00010000100111" => data_out <= "100";
            when "00010000101000" => data_out <= "100";
            when "00010000101001" => data_out <= "100";
            when "00010000101010" => data_out <= "000";
            when "00010000101011" => data_out <= "000";
            when "00010000101100" => data_out <= "000";
            when "00010000101101" => data_out <= "000";
            when "00010000101110" => data_out <= "000";
            when "00010000101111" => data_out <= "000";
            when "00010000110000" => data_out <= "100";
            when "00010000110001" => data_out <= "100";
            when "00010000110010" => data_out <= "111";
            when "00010000110011" => data_out <= "111";
            when "00010000110100" => data_out <= "111";
            when "00010000110101" => data_out <= "111";
            when "00010000110110" => data_out <= "111";
            when "00010000110111" => data_out <= "111";
            when "00010000111000" => data_out <= "111";
            when "00010000111001" => data_out <= "111";
            when "00010000111010" => data_out <= "111";
            when "00010000111011" => data_out <= "111";
            when "00010000111100" => data_out <= "111";
            when "00010000111101" => data_out <= "111";
            when "00010000111110" => data_out <= "111";
            when "00010000111111" => data_out <= "111";
            when "00010001000000" => data_out <= "111";
            when "00010001000001" => data_out <= "111";
            when "00010001000010" => data_out <= "111";
            when "00010001000011" => data_out <= "111";
            when "00010001000100" => data_out <= "111";
            when "00010001000101" => data_out <= "111";
            when "00010001000110" => data_out <= "111";
            when "00010001000111" => data_out <= "111";
            when "00010001001000" => data_out <= "000";
            when "00010001001001" => data_out <= "000";
            when "00010001001010" => data_out <= "000";
            when "00010001001011" => data_out <= "000";
            when "00010001001100" => data_out <= "000";
            when "00010001001101" => data_out <= "000";
            when "00010001001110" => data_out <= "000";
            when "00010001001111" => data_out <= "000";
            when "00010001010000" => data_out <= "000";
            when "00010001010001" => data_out <= "000";
            when "00010001010010" => data_out <= "000";
            when "00010001010011" => data_out <= "000";
            when "00010001010100" => data_out <= "000";
            when "00010001010101" => data_out <= "000";
            when "00010001010110" => data_out <= "000";
            when "00010001010111" => data_out <= "000";
            when "00010001011000" => data_out <= "000";
            when "00010001011001" => data_out <= "000";
            when "00010001011010" => data_out <= "000";
            when "00010001011011" => data_out <= "000";
            when "00010001011100" => data_out <= "000";
            when "00010001011101" => data_out <= "000";
            when "00010001011110" => data_out <= "000";
            when "00010001011111" => data_out <= "000";
            when "00010001100000" => data_out <= "000";
            when "00010001100001" => data_out <= "000";
            when "00010001100010" => data_out <= "000";
            when "00010001100011" => data_out <= "000";
            when "00010001100100" => data_out <= "000";
            when "00010001100101" => data_out <= "000";
            when "00010001100110" => data_out <= "000";
            when "00010001100111" => data_out <= "000";
            when "00010001101000" => data_out <= "000";
            when "00010001101001" => data_out <= "000";
            when "00010001101010" => data_out <= "000";
            when "00010001101011" => data_out <= "000";
            when "00010001101100" => data_out <= "000";
            when "00010001101101" => data_out <= "000";
            when "00010001101110" => data_out <= "000";
            when "00010001101111" => data_out <= "000";
            when "00010001110000" => data_out <= "000";
            when "00010001110001" => data_out <= "000";
            when "00010001110010" => data_out <= "000";
            when "00010001110011" => data_out <= "000";
            when "00010001110100" => data_out <= "000";
            when "00010001110101" => data_out <= "000";
            when "00010001110110" => data_out <= "000";
            when "00010001110111" => data_out <= "000";
            when "00010001111000" => data_out <= "000";
            when "00010001111001" => data_out <= "000";
            when "00010001111010" => data_out <= "000";
            when "00010001111011" => data_out <= "000";
            when "00010001111100" => data_out <= "000";
            when "00010001111101" => data_out <= "000";
            when "00010001111110" => data_out <= "000";
            when "00010001111111" => data_out <= "000";
            when "00010010000000" => data_out <= "000";
            when "00010010000001" => data_out <= "000";
            when "00010010000010" => data_out <= "000";
            when "00010010000011" => data_out <= "000";
            when "00010010000100" => data_out <= "000";
            when "00010010000101" => data_out <= "000";
            when "00010010000110" => data_out <= "000";
            when "00010010000111" => data_out <= "000";
            when "00010010001000" => data_out <= "000";
            when "00010010001001" => data_out <= "000";
            when "00010010001010" => data_out <= "000";
            when "00010010001011" => data_out <= "000";
            when "00010010001100" => data_out <= "000";
            when "00010010001101" => data_out <= "000";
            when "00010010001110" => data_out <= "000";
            when "00010010001111" => data_out <= "111";
            when "00010010010000" => data_out <= "111";
            when "00010010010001" => data_out <= "111";
            when "00010010010010" => data_out <= "111";
            when "00010010010011" => data_out <= "111";
            when "00010010010100" => data_out <= "111";
            when "00010010010101" => data_out <= "111";
            when "00010010010110" => data_out <= "111";
            when "00010010010111" => data_out <= "100";
            when "00010010011000" => data_out <= "100";
            when "00010010011001" => data_out <= "100";
            when "00010010011010" => data_out <= "100";
            when "00010010011011" => data_out <= "100";
            when "00010010011100" => data_out <= "100";
            when "00010010011101" => data_out <= "100";
            when "00010010011110" => data_out <= "100";
            when "00010010011111" => data_out <= "100";
            when "00010010100000" => data_out <= "100";
            when "00010010100001" => data_out <= "100";
            when "00010010100010" => data_out <= "100";
            when "00010010100011" => data_out <= "100";
            when "00010010100100" => data_out <= "100";
            when "00010010100101" => data_out <= "100";
            when "00010010100110" => data_out <= "100";
            when "00010010100111" => data_out <= "100";
            when "00010010101000" => data_out <= "100";
            when "00010010101001" => data_out <= "100";
            when "00010010101010" => data_out <= "100";
            when "00010010101011" => data_out <= "100";
            when "00010010101100" => data_out <= "100";
            when "00010010101101" => data_out <= "100";
            when "00010010101110" => data_out <= "100";
            when "00010010101111" => data_out <= "100";
            when "00010010110000" => data_out <= "100";
            when "00010010110001" => data_out <= "100";
            when "00010010110010" => data_out <= "100";
            when "00010010110011" => data_out <= "100";
            when "00010010110100" => data_out <= "100";
            when "00010010110101" => data_out <= "100";
            when "00010010110110" => data_out <= "111";
            when "00010010110111" => data_out <= "111";
            when "00010010111000" => data_out <= "111";
            when "00010010111001" => data_out <= "111";
            when "00010010111010" => data_out <= "111";
            when "00010010111011" => data_out <= "111";
            when "00010010111100" => data_out <= "111";
            when "00010010111101" => data_out <= "111";
            when "00010010111110" => data_out <= "111";
            when "00010010111111" => data_out <= "000";
            when "00010011000000" => data_out <= "000";
            when "00010011000001" => data_out <= "000";
            when "00010011000010" => data_out <= "000";
            when "00010011000011" => data_out <= "000";
            when "00010011000100" => data_out <= "000";
            when "00010011000101" => data_out <= "000";
            when "00010011000110" => data_out <= "000";
            when "00010011000111" => data_out <= "000";
            when "00010011001000" => data_out <= "000";
            when "00010011001001" => data_out <= "000";
            when "00010011001010" => data_out <= "000";
            when "00010011001011" => data_out <= "000";
            when "00010011001100" => data_out <= "000";
            when "00010011001101" => data_out <= "000";
            when "00010011001110" => data_out <= "111";
            when "00010011001111" => data_out <= "000";
            when "00010011010000" => data_out <= "000";
            when "00010011010001" => data_out <= "000";
            when "00010011010010" => data_out <= "000";
            when "00010011010011" => data_out <= "000";
            when "00010011010100" => data_out <= "000";
            when "00010011010101" => data_out <= "000";
            when "00010011010110" => data_out <= "000";
            when "00010011010111" => data_out <= "000";
            when "00010011011000" => data_out <= "000";
            when "00010011011001" => data_out <= "000";
            when "00010011011010" => data_out <= "000";
            when "00010011011011" => data_out <= "000";
            when "00010011011100" => data_out <= "000";
            when "00010011011101" => data_out <= "000";
            when "00010011011110" => data_out <= "000";
            when "00010011011111" => data_out <= "000";
            when "00010011100000" => data_out <= "000";
            when "00010011100001" => data_out <= "000";
            when "00010011100010" => data_out <= "000";
            when "00010011100011" => data_out <= "000";
            when "00010011100100" => data_out <= "000";
            when "00010011100101" => data_out <= "000";
            when "00010011100110" => data_out <= "000";
            when "00010011100111" => data_out <= "000";
            when "00010011101000" => data_out <= "000";
            when "00010011101001" => data_out <= "000";
            when "00010011101010" => data_out <= "000";
            when "00010011101011" => data_out <= "000";
            when "00010011101100" => data_out <= "000";
            when "00010011101101" => data_out <= "000";
            when "00010011101110" => data_out <= "000";
            when "00010011101111" => data_out <= "000";
            when "00010011110000" => data_out <= "000";
            when "00010011110001" => data_out <= "000";
            when "00010011110010" => data_out <= "000";
            when "00010011110011" => data_out <= "000";
            when "00010011110100" => data_out <= "000";
            when "00010011110101" => data_out <= "000";
            when "00010011110110" => data_out <= "000";
            when "00010011110111" => data_out <= "000";
            when "00010011111000" => data_out <= "000";
            when "00010011111001" => data_out <= "000";
            when "00010011111010" => data_out <= "000";
            when "00010011111011" => data_out <= "000";
            when "00010011111100" => data_out <= "000";
            when "00010011111101" => data_out <= "000";
            when "00010011111110" => data_out <= "000";
            when "00010011111111" => data_out <= "000";
            when "00010100000000" => data_out <= "000";
            when "00010100000001" => data_out <= "000";
            when "00010100000010" => data_out <= "000";
            when "00010100000011" => data_out <= "000";
            when "00010100000100" => data_out <= "000";
            when "00010100000101" => data_out <= "000";
            when "00010100000110" => data_out <= "000";
            when "00010100000111" => data_out <= "000";
            when "00010100001000" => data_out <= "000";
            when "00010100001001" => data_out <= "000";
            when "00010100001010" => data_out <= "000";
            when "00010100001011" => data_out <= "000";
            when "00010100001100" => data_out <= "000";
            when "00010100001101" => data_out <= "000";
            when "00010100001110" => data_out <= "000";
            when "00010100001111" => data_out <= "000";
            when "00010100010000" => data_out <= "000";
            when "00010100010001" => data_out <= "000";
            when "00010100010010" => data_out <= "000";
            when "00010100010011" => data_out <= "000";
            when "00010100010100" => data_out <= "000";
            when "00010100010101" => data_out <= "000";
            when "00010100010110" => data_out <= "000";
            when "00010100010111" => data_out <= "111";
            when "00010100011000" => data_out <= "111";
            when "00010100011001" => data_out <= "111";
            when "00010100011010" => data_out <= "111";
            when "00010100011011" => data_out <= "111";
            when "00010100011100" => data_out <= "111";
            when "00010100011101" => data_out <= "111";
            when "00010100011110" => data_out <= "111";
            when "00010100011111" => data_out <= "111";
            when "00010100100000" => data_out <= "100";
            when "00010100100001" => data_out <= "100";
            when "00010100100010" => data_out <= "100";
            when "00010100100011" => data_out <= "100";
            when "00010100100100" => data_out <= "100";
            when "00010100100101" => data_out <= "100";
            when "00010100100110" => data_out <= "100";
            when "00010100100111" => data_out <= "100";
            when "00010100101000" => data_out <= "100";
            when "00010100101001" => data_out <= "100";
            when "00010100101010" => data_out <= "100";
            when "00010100101011" => data_out <= "100";
            when "00010100101100" => data_out <= "100";
            when "00010100101101" => data_out <= "100";
            when "00010100101110" => data_out <= "100";
            when "00010100101111" => data_out <= "100";
            when "00010100110000" => data_out <= "100";
            when "00010100110001" => data_out <= "100";
            when "00010100110010" => data_out <= "111";
            when "00010100110011" => data_out <= "111";
            when "00010100110100" => data_out <= "111";
            when "00010100110101" => data_out <= "111";
            when "00010100110110" => data_out <= "111";
            when "00010100110111" => data_out <= "111";
            when "00010100111000" => data_out <= "111";
            when "00010100111001" => data_out <= "111";
            when "00010100111010" => data_out <= "111";
            when "00010100111011" => data_out <= "000";
            when "00010100111100" => data_out <= "000";
            when "00010100111101" => data_out <= "000";
            when "00010100111110" => data_out <= "000";
            when "00010100111111" => data_out <= "000";
            when "00010101000000" => data_out <= "000";
            when "00010101000001" => data_out <= "000";
            when "00010101000010" => data_out <= "000";
            when "00010101000011" => data_out <= "000";
            when "00010101000100" => data_out <= "000";
            when "00010101000101" => data_out <= "000";
            when "00010101000110" => data_out <= "000";
            when "00010101000111" => data_out <= "000";
            when "00010101001000" => data_out <= "000";
            when "00010101001001" => data_out <= "000";
            when "00010101001010" => data_out <= "000";
            when "00010101001011" => data_out <= "000";
            when "00010101001100" => data_out <= "000";
            when "00010101001101" => data_out <= "000";
            when "00010101001110" => data_out <= "111";
            when "00010101001111" => data_out <= "111";
            when "00010101010000" => data_out <= "000";
            when "00010101010001" => data_out <= "111";
            when "00010101010010" => data_out <= "000";
            when "00010101010011" => data_out <= "000";
            when "00010101010100" => data_out <= "000";
            when "00010101010101" => data_out <= "000";
            when "00010101010110" => data_out <= "000";
            when "00010101010111" => data_out <= "000";
            when "00010101011000" => data_out <= "000";
            when "00010101011001" => data_out <= "000";
            when "00010101011010" => data_out <= "000";
            when "00010101011011" => data_out <= "000";
            when "00010101011100" => data_out <= "000";
            when "00010101011101" => data_out <= "000";
            when "00010101011110" => data_out <= "000";
            when "00010101011111" => data_out <= "000";
            when "00010101100000" => data_out <= "000";
            when "00010101100001" => data_out <= "000";
            when "00010101100010" => data_out <= "000";
            when "00010101100011" => data_out <= "000";
            when "00010101100100" => data_out <= "000";
            when "00010101100101" => data_out <= "000";
            when "00010101100110" => data_out <= "000";
            when "00010101100111" => data_out <= "000";
            when "00010101101000" => data_out <= "000";
            when "00010101101001" => data_out <= "000";
            when "00010101101010" => data_out <= "000";
            when "00010101101011" => data_out <= "000";
            when "00010101101100" => data_out <= "000";
            when "00010101101101" => data_out <= "000";
            when "00010101101110" => data_out <= "000";
            when "00010101101111" => data_out <= "000";
            when "00010101110000" => data_out <= "000";
            when "00010101110001" => data_out <= "000";
            when "00010101110010" => data_out <= "000";
            when "00010101110011" => data_out <= "000";
            when "00010101110100" => data_out <= "000";
            when "00010101110101" => data_out <= "000";
            when "00010101110110" => data_out <= "000";
            when "00010101110111" => data_out <= "000";
            when "00010101111000" => data_out <= "000";
            when "00010101111001" => data_out <= "000";
            when "00010101111010" => data_out <= "000";
            when "00010101111011" => data_out <= "000";
            when "00010101111100" => data_out <= "000";
            when "00010101111101" => data_out <= "000";
            when "00010101111110" => data_out <= "000";
            when "00010101111111" => data_out <= "000";
            when "00010110000000" => data_out <= "000";
            when "00010110000001" => data_out <= "000";
            when "00010110000010" => data_out <= "000";
            when "00010110000011" => data_out <= "000";
            when "00010110000100" => data_out <= "000";
            when "00010110000101" => data_out <= "000";
            when "00010110000110" => data_out <= "000";
            when "00010110000111" => data_out <= "000";
            when "00010110001000" => data_out <= "000";
            when "00010110001001" => data_out <= "000";
            when "00010110001010" => data_out <= "000";
            when "00010110001011" => data_out <= "000";
            when "00010110001100" => data_out <= "000";
            when "00010110001101" => data_out <= "000";
            when "00010110001110" => data_out <= "000";
            when "00010110001111" => data_out <= "000";
            when "00010110010000" => data_out <= "000";
            when "00010110010001" => data_out <= "000";
            when "00010110010010" => data_out <= "000";
            when "00010110010011" => data_out <= "000";
            when "00010110010100" => data_out <= "000";
            when "00010110010101" => data_out <= "000";
            when "00010110010110" => data_out <= "000";
            when "00010110010111" => data_out <= "000";
            when "00010110011000" => data_out <= "000";
            when "00010110011001" => data_out <= "000";
            when "00010110011010" => data_out <= "000";
            when "00010110011011" => data_out <= "000";
            when "00010110011100" => data_out <= "000";
            when "00010110011101" => data_out <= "000";
            when "00010110011110" => data_out <= "000";
            when "00010110011111" => data_out <= "000";
            when "00010110100000" => data_out <= "111";
            when "00010110100001" => data_out <= "111";
            when "00010110100010" => data_out <= "111";
            when "00010110100011" => data_out <= "111";
            when "00010110100100" => data_out <= "111";
            when "00010110100101" => data_out <= "111";
            when "00010110100110" => data_out <= "111";
            when "00010110100111" => data_out <= "111";
            when "00010110101000" => data_out <= "111";
            when "00010110101001" => data_out <= "111";
            when "00010110101010" => data_out <= "111";
            when "00010110101011" => data_out <= "111";
            when "00010110101100" => data_out <= "111";
            when "00010110101101" => data_out <= "111";
            when "00010110101110" => data_out <= "111";
            when "00010110101111" => data_out <= "111";
            when "00010110110000" => data_out <= "111";
            when "00010110110001" => data_out <= "111";
            when "00010110110010" => data_out <= "000";
            when "00010110110011" => data_out <= "000";
            when "00010110110100" => data_out <= "000";
            when "00010110110101" => data_out <= "000";
            when "00010110110110" => data_out <= "000";
            when "00010110110111" => data_out <= "000";
            when "00010110111000" => data_out <= "000";
            when "00010110111001" => data_out <= "000";
            when "00010110111010" => data_out <= "000";
            when "00010110111011" => data_out <= "000";
            when "00010110111100" => data_out <= "000";
            when "00010110111101" => data_out <= "000";
            when "00010110111110" => data_out <= "000";
            when "00010110111111" => data_out <= "000";
            when "00010111000000" => data_out <= "000";
            when "00010111000001" => data_out <= "000";
            when "00010111000010" => data_out <= "000";
            when "00010111000011" => data_out <= "000";
            when "00010111000100" => data_out <= "000";
            when "00010111000101" => data_out <= "000";
            when "00010111000110" => data_out <= "000";
            when "00010111000111" => data_out <= "000";
            when "00010111001000" => data_out <= "000";
            when "00010111001001" => data_out <= "000";
            when "00010111001010" => data_out <= "000";
            when "00010111001011" => data_out <= "000";
            when "00010111001100" => data_out <= "000";
            when "00010111001101" => data_out <= "000";
            when "00010111001110" => data_out <= "111";
            when "00010111001111" => data_out <= "000";
            when "00010111010000" => data_out <= "000";
            when "00010111010001" => data_out <= "000";
            when "00010111010010" => data_out <= "111";
            when "00010111010011" => data_out <= "111";
            when "00010111010100" => data_out <= "000";
            when "00010111010101" => data_out <= "000";
            when "00010111010110" => data_out <= "000";
            when "00010111010111" => data_out <= "000";
            when "00010111011000" => data_out <= "000";
            when "00010111011001" => data_out <= "000";
            when "00010111011010" => data_out <= "000";
            when "00010111011011" => data_out <= "000";
            when "00010111011100" => data_out <= "000";
            when "00010111011101" => data_out <= "000";
            when "00010111011110" => data_out <= "000";
            when "00010111011111" => data_out <= "000";
            when "00010111100000" => data_out <= "000";
            when "00010111100001" => data_out <= "000";
            when "00010111100010" => data_out <= "000";
            when "00010111100011" => data_out <= "000";
            when "00010111100100" => data_out <= "000";
            when "00010111100101" => data_out <= "000";
            when "00010111100110" => data_out <= "000";
            when "00010111100111" => data_out <= "000";
            when "00010111101000" => data_out <= "000";
            when "00010111101001" => data_out <= "000";
            when "00010111101010" => data_out <= "000";
            when "00010111101011" => data_out <= "000";
            when "00010111101100" => data_out <= "000";
            when "00010111101101" => data_out <= "000";
            when "00010111101110" => data_out <= "000";
            when "00010111101111" => data_out <= "000";
            when "00010111110000" => data_out <= "000";
            when "00010111110001" => data_out <= "000";
            when "00010111110010" => data_out <= "000";
            when "00010111110011" => data_out <= "000";
            when "00010111110100" => data_out <= "000";
            when "00010111110101" => data_out <= "000";
            when "00010111110110" => data_out <= "000";
            when "00010111110111" => data_out <= "000";
            when "00010111111000" => data_out <= "000";
            when "00010111111001" => data_out <= "000";
            when "00010111111010" => data_out <= "000";
            when "00010111111011" => data_out <= "000";
            when "00010111111100" => data_out <= "000";
            when "00010111111101" => data_out <= "000";
            when "00010111111110" => data_out <= "000";
            when "00010111111111" => data_out <= "000";
            when "00011000000000" => data_out <= "000";
            when "00011000000001" => data_out <= "000";
            when "00011000000010" => data_out <= "000";
            when "00011000000011" => data_out <= "000";
            when "00011000000100" => data_out <= "000";
            when "00011000000101" => data_out <= "000";
            when "00011000000110" => data_out <= "000";
            when "00011000000111" => data_out <= "000";
            when "00011000001000" => data_out <= "000";
            when "00011000001001" => data_out <= "000";
            when "00011000001010" => data_out <= "000";
            when "00011000001011" => data_out <= "000";
            when "00011000001100" => data_out <= "000";
            when "00011000001101" => data_out <= "000";
            when "00011000001110" => data_out <= "000";
            when "00011000001111" => data_out <= "000";
            when "00011000010000" => data_out <= "000";
            when "00011000010001" => data_out <= "000";
            when "00011000010010" => data_out <= "000";
            when "00011000010011" => data_out <= "000";
            when "00011000010100" => data_out <= "000";
            when "00011000010101" => data_out <= "000";
            when "00011000010110" => data_out <= "000";
            when "00011000010111" => data_out <= "000";
            when "00011000011000" => data_out <= "000";
            when "00011000011001" => data_out <= "000";
            when "00011000011010" => data_out <= "000";
            when "00011000011011" => data_out <= "000";
            when "00011000011100" => data_out <= "000";
            when "00011000011101" => data_out <= "000";
            when "00011000011110" => data_out <= "000";
            when "00011000011111" => data_out <= "000";
            when "00011000100000" => data_out <= "000";
            when "00011000100001" => data_out <= "000";
            when "00011000100010" => data_out <= "000";
            when "00011000100011" => data_out <= "000";
            when "00011000100100" => data_out <= "000";
            when "00011000100101" => data_out <= "000";
            when "00011000100110" => data_out <= "000";
            when "00011000100111" => data_out <= "000";
            when "00011000101000" => data_out <= "000";
            when "00011000101001" => data_out <= "000";
            when "00011000101010" => data_out <= "000";
            when "00011000101011" => data_out <= "000";
            when "00011000101100" => data_out <= "000";
            when "00011000101101" => data_out <= "000";
            when "00011000101110" => data_out <= "000";
            when "00011000101111" => data_out <= "000";
            when "00011000110000" => data_out <= "000";
            when "00011000110001" => data_out <= "000";
            when "00011000110010" => data_out <= "000";
            when "00011000110011" => data_out <= "000";
            when "00011000110100" => data_out <= "000";
            when "00011000110101" => data_out <= "000";
            when "00011000110110" => data_out <= "000";
            when "00011000110111" => data_out <= "000";
            when "00011000111000" => data_out <= "000";
            when "00011000111001" => data_out <= "000";
            when "00011000111010" => data_out <= "000";
            when "00011000111011" => data_out <= "000";
            when "00011000111100" => data_out <= "000";
            when "00011000111101" => data_out <= "000";
            when "00011000111110" => data_out <= "000";
            when "00011000111111" => data_out <= "000";
            when "00011001000000" => data_out <= "000";
            when "00011001000001" => data_out <= "000";
            when "00011001000010" => data_out <= "000";
            when "00011001000011" => data_out <= "000";
            when "00011001000100" => data_out <= "000";
            when "00011001000101" => data_out <= "000";
            when "00011001000110" => data_out <= "000";
            when "00011001000111" => data_out <= "000";
            when "00011001001000" => data_out <= "000";
            when "00011001001001" => data_out <= "000";
            when "00011001001010" => data_out <= "000";
            when "00011001001011" => data_out <= "000";
            when "00011001001100" => data_out <= "000";
            when "00011001001101" => data_out <= "000";
            when "00011001001110" => data_out <= "111";
            when "00011001001111" => data_out <= "000";
            when "00011001010000" => data_out <= "000";
            when "00011001010001" => data_out <= "000";
            when "00011001010010" => data_out <= "000";
            when "00011001010011" => data_out <= "000";
            when "00011001010100" => data_out <= "000";
            when "00011001010101" => data_out <= "000";
            when "00011001010110" => data_out <= "000";
            when "00011001010111" => data_out <= "000";
            when "00011001011000" => data_out <= "000";
            when "00011001011001" => data_out <= "000";
            when "00011001011010" => data_out <= "000";
            when "00011001011011" => data_out <= "000";
            when "00011001011100" => data_out <= "000";
            when "00011001011101" => data_out <= "000";
            when "00011001011110" => data_out <= "000";
            when "00011001011111" => data_out <= "000";
            when "00011001100000" => data_out <= "000";
            when "00011001100001" => data_out <= "000";
            when "00011001100010" => data_out <= "000";
            when "00011001100011" => data_out <= "000";
            when "00011001100100" => data_out <= "000";
            when "00011001100101" => data_out <= "000";
            when "00011001100110" => data_out <= "000";
            when "00011001100111" => data_out <= "000";
            when "00011001101000" => data_out <= "000";
            when "00011001101001" => data_out <= "000";
            when "00011001101010" => data_out <= "000";
            when "00011001101011" => data_out <= "000";
            when "00011001101100" => data_out <= "000";
            when "00011001101101" => data_out <= "000";
            when "00011001101110" => data_out <= "000";
            when "00011001101111" => data_out <= "000";
            when "00011001110000" => data_out <= "000";
            when "00011001110001" => data_out <= "000";
            when "00011001110010" => data_out <= "000";
            when "00011001110011" => data_out <= "000";
            when "00011001110100" => data_out <= "000";
            when "00011001110101" => data_out <= "000";
            when "00011001110110" => data_out <= "000";
            when "00011001110111" => data_out <= "000";
            when "00011001111000" => data_out <= "000";
            when "00011001111001" => data_out <= "000";
            when "00011001111010" => data_out <= "000";
            when "00011001111011" => data_out <= "000";
            when "00011001111100" => data_out <= "000";
            when "00011001111101" => data_out <= "000";
            when "00011001111110" => data_out <= "000";
            when "00011001111111" => data_out <= "000";
            when "00011010000000" => data_out <= "000";
            when "00011010000001" => data_out <= "000";
            when "00011010000010" => data_out <= "000";
            when "00011010000011" => data_out <= "000";
            when "00011010000100" => data_out <= "000";
            when "00011010000101" => data_out <= "000";
            when "00011010000110" => data_out <= "000";
            when "00011010000111" => data_out <= "000";
            when "00011010001000" => data_out <= "000";
            when "00011010001001" => data_out <= "000";
            when "00011010001010" => data_out <= "000";
            when "00011010001011" => data_out <= "000";
            when "00011010001100" => data_out <= "000";
            when "00011010001101" => data_out <= "000";
            when "00011010001110" => data_out <= "000";
            when "00011010001111" => data_out <= "000";
            when "00011010010000" => data_out <= "000";
            when "00011010010001" => data_out <= "000";
            when "00011010010010" => data_out <= "000";
            when "00011010010011" => data_out <= "000";
            when "00011010010100" => data_out <= "000";
            when "00011010010101" => data_out <= "000";
            when "00011010010110" => data_out <= "000";
            when "00011010010111" => data_out <= "000";
            when "00011010011000" => data_out <= "000";
            when "00011010011001" => data_out <= "000";
            when "00011010011010" => data_out <= "000";
            when "00011010011011" => data_out <= "000";
            when "00011010011100" => data_out <= "000";
            when "00011010011101" => data_out <= "000";
            when "00011010011110" => data_out <= "000";
            when "00011010011111" => data_out <= "000";
            when "00011010100000" => data_out <= "000";
            when "00011010100001" => data_out <= "000";
            when "00011010100010" => data_out <= "000";
            when "00011010100011" => data_out <= "000";
            when "00011010100100" => data_out <= "000";
            when "00011010100101" => data_out <= "000";
            when "00011010100110" => data_out <= "000";
            when "00011010100111" => data_out <= "000";
            when "00011010101000" => data_out <= "000";
            when "00011010101001" => data_out <= "000";
            when "00011010101010" => data_out <= "000";
            when "00011010101011" => data_out <= "000";
            when "00011010101100" => data_out <= "000";
            when "00011010101101" => data_out <= "000";
            when "00011010101110" => data_out <= "000";
            when "00011010101111" => data_out <= "000";
            when "00011010110000" => data_out <= "000";
            when "00011010110001" => data_out <= "000";
            when "00011010110010" => data_out <= "000";
            when "00011010110011" => data_out <= "000";
            when "00011010110100" => data_out <= "000";
            when "00011010110101" => data_out <= "000";
            when "00011010110110" => data_out <= "000";
            when "00011010110111" => data_out <= "000";
            when "00011010111000" => data_out <= "000";
            when "00011010111001" => data_out <= "000";
            when "00011010111010" => data_out <= "000";
            when "00011010111011" => data_out <= "000";
            when "00011010111100" => data_out <= "000";
            when "00011010111101" => data_out <= "000";
            when "00011010111110" => data_out <= "000";
            when "00011010111111" => data_out <= "000";
            when "00011011000000" => data_out <= "000";
            when "00011011000001" => data_out <= "000";
            when "00011011000010" => data_out <= "000";
            when "00011011000011" => data_out <= "000";
            when "00011011000100" => data_out <= "000";
            when "00011011000101" => data_out <= "000";
            when "00011011000110" => data_out <= "000";
            when "00011011000111" => data_out <= "000";
            when "00011011001000" => data_out <= "000";
            when "00011011001001" => data_out <= "000";
            when "00011011001010" => data_out <= "000";
            when "00011011001011" => data_out <= "000";
            when "00011011001100" => data_out <= "000";
            when "00011011001101" => data_out <= "000";
            when "00011011001110" => data_out <= "000";
            when "00011011001111" => data_out <= "000";
            when "00011011010000" => data_out <= "000";
            when "00011011010001" => data_out <= "000";
            when "00011011010010" => data_out <= "000";
            when "00011011010011" => data_out <= "000";
            when "00011011010100" => data_out <= "000";
            when "00011011010101" => data_out <= "000";
            when "00011011010110" => data_out <= "000";
            when "00011011010111" => data_out <= "000";
            when "00011011011000" => data_out <= "000";
            when "00011011011001" => data_out <= "000";
            when "00011011011010" => data_out <= "000";
            when "00011011011011" => data_out <= "000";
            when "00011011011100" => data_out <= "000";
            when "00011011011101" => data_out <= "000";
            when "00011011011110" => data_out <= "000";
            when "00011011011111" => data_out <= "000";
            when "00011011100000" => data_out <= "000";
            when "00011011100001" => data_out <= "000";
            when "00011011100010" => data_out <= "000";
            when "00011011100011" => data_out <= "000";
            when "00011011100100" => data_out <= "000";
            when "00011011100101" => data_out <= "000";
            when "00011011100110" => data_out <= "000";
            when "00011011100111" => data_out <= "000";
            when "00011011101000" => data_out <= "000";
            when "00011011101001" => data_out <= "000";
            when "00011011101010" => data_out <= "000";
            when "00011011101011" => data_out <= "000";
            when "00011011101100" => data_out <= "000";
            when "00011011101101" => data_out <= "000";
            when "00011011101110" => data_out <= "000";
            when "00011011101111" => data_out <= "000";
            when "00011011110000" => data_out <= "000";
            when "00011011110001" => data_out <= "000";
            when "00011011110010" => data_out <= "000";
            when "00011011110011" => data_out <= "000";
            when "00011011110100" => data_out <= "000";
            when "00011011110101" => data_out <= "000";
            when "00011011110110" => data_out <= "000";
            when "00011011110111" => data_out <= "000";
            when "00011011111000" => data_out <= "000";
            when "00011011111001" => data_out <= "000";
            when "00011011111010" => data_out <= "000";
            when "00011011111011" => data_out <= "000";
            when "00011011111100" => data_out <= "000";
            when "00011011111101" => data_out <= "000";
            when "00011011111110" => data_out <= "000";
            when "00011011111111" => data_out <= "000";
            when "00011100000000" => data_out <= "000";
            when "00011100000001" => data_out <= "000";
            when "00011100000010" => data_out <= "000";
            when "00011100000011" => data_out <= "000";
            when "00011100000100" => data_out <= "000";
            when "00011100000101" => data_out <= "000";
            when "00011100000110" => data_out <= "000";
            when "00011100000111" => data_out <= "000";
            when "00011100001000" => data_out <= "000";
            when "00011100001001" => data_out <= "000";
            when "00011100001010" => data_out <= "000";
            when "00011100001011" => data_out <= "000";
            when "00011100001100" => data_out <= "000";
            when "00011100001101" => data_out <= "000";
            when "00011100001110" => data_out <= "000";
            when "00011100001111" => data_out <= "000";
            when "00011100010000" => data_out <= "000";
            when "00011100010001" => data_out <= "000";
            when "00011100010010" => data_out <= "000";
            when "00011100010011" => data_out <= "000";
            when "00011100010100" => data_out <= "000";
            when "00011100010101" => data_out <= "000";
            when "00011100010110" => data_out <= "000";
            when "00011100010111" => data_out <= "000";
            when "00011100011000" => data_out <= "000";
            when "00011100011001" => data_out <= "000";
            when "00011100011010" => data_out <= "000";
            when "00011100011011" => data_out <= "000";
            when "00011100011100" => data_out <= "000";
            when "00011100011101" => data_out <= "000";
            when "00011100011110" => data_out <= "000";
            when "00011100011111" => data_out <= "000";
            when "00011100100000" => data_out <= "000";
            when "00011100100001" => data_out <= "000";
            when "00011100100010" => data_out <= "000";
            when "00011100100011" => data_out <= "000";
            when "00011100100100" => data_out <= "000";
            when "00011100100101" => data_out <= "000";
            when "00011100100110" => data_out <= "000";
            when "00011100100111" => data_out <= "000";
            when "00011100101000" => data_out <= "000";
            when "00011100101001" => data_out <= "000";
            when "00011100101010" => data_out <= "000";
            when "00011100101011" => data_out <= "000";
            when "00011100101100" => data_out <= "000";
            when "00011100101101" => data_out <= "000";
            when "00011100101110" => data_out <= "000";
            when "00011100101111" => data_out <= "000";
            when "00011100110000" => data_out <= "000";
            when "00011100110001" => data_out <= "000";
            when "00011100110010" => data_out <= "000";
            when "00011100110011" => data_out <= "000";
            when "00011100110100" => data_out <= "000";
            when "00011100110101" => data_out <= "000";
            when "00011100110110" => data_out <= "000";
            when "00011100110111" => data_out <= "000";
            when "00011100111000" => data_out <= "000";
            when "00011100111001" => data_out <= "000";
            when "00011100111010" => data_out <= "000";
            when "00011100111011" => data_out <= "000";
            when "00011100111100" => data_out <= "000";
            when "00011100111101" => data_out <= "000";
            when "00011100111110" => data_out <= "000";
            when "00011100111111" => data_out <= "000";
            when "00011101000000" => data_out <= "000";
            when "00011101000001" => data_out <= "000";
            when "00011101000010" => data_out <= "000";
            when "00011101000011" => data_out <= "000";
            when "00011101000100" => data_out <= "000";
            when "00011101000101" => data_out <= "000";
            when "00011101000110" => data_out <= "000";
            when "00011101000111" => data_out <= "000";
            when "00011101001000" => data_out <= "000";
            when "00011101001001" => data_out <= "000";
            when "00011101001010" => data_out <= "000";
            when "00011101001011" => data_out <= "000";
            when "00011101001100" => data_out <= "000";
            when "00011101001101" => data_out <= "000";
            when "00011101001110" => data_out <= "000";
            when "00011101001111" => data_out <= "000";
            when "00011101010000" => data_out <= "000";
            when "00011101010001" => data_out <= "000";
            when "00011101010010" => data_out <= "000";
            when "00011101010011" => data_out <= "000";
            when "00011101010100" => data_out <= "000";
            when "00011101010101" => data_out <= "000";
            when "00011101010110" => data_out <= "000";
            when "00011101010111" => data_out <= "000";
            when "00011101011000" => data_out <= "000";
            when "00011101011001" => data_out <= "000";
            when "00011101011010" => data_out <= "000";
            when "00011101011011" => data_out <= "000";
            when "00011101011100" => data_out <= "000";
            when "00011101011101" => data_out <= "000";
            when "00011101011110" => data_out <= "000";
            when "00011101011111" => data_out <= "000";
            when "00011101100000" => data_out <= "000";
            when "00011101100001" => data_out <= "000";
            when "00011101100010" => data_out <= "000";
            when "00011101100011" => data_out <= "000";
            when "00011101100100" => data_out <= "000";
            when "00011101100101" => data_out <= "000";
            when "00011101100110" => data_out <= "000";
            when "00011101100111" => data_out <= "000";
            when "00011101101000" => data_out <= "000";
            when "00011101101001" => data_out <= "000";
            when "00011101101010" => data_out <= "000";
            when "00011101101011" => data_out <= "000";
            when "00011101101100" => data_out <= "000";
            when "00011101101101" => data_out <= "000";
            when "00011101101110" => data_out <= "000";
            when "00011101101111" => data_out <= "000";
            when "00011101110000" => data_out <= "000";
            when "00011101110001" => data_out <= "000";
            when "00011101110010" => data_out <= "000";
            when "00011101110011" => data_out <= "000";
            when "00011101110100" => data_out <= "000";
            when "00011101110101" => data_out <= "000";
            when "00011101110110" => data_out <= "000";
            when "00011101110111" => data_out <= "000";
            when "00011101111000" => data_out <= "000";
            when "00011101111001" => data_out <= "000";
            when "00011101111010" => data_out <= "000";
            when "00011101111011" => data_out <= "000";
            when "00011101111100" => data_out <= "000";
            when "00011101111101" => data_out <= "000";
            when "00011101111110" => data_out <= "000";
            when "00011101111111" => data_out <= "000";
            when "00011110000000" => data_out <= "000";
            when "00011110000001" => data_out <= "000";
            when "00011110000010" => data_out <= "000";
            when "00011110000011" => data_out <= "000";
            when "00011110000100" => data_out <= "000";
            when "00011110000101" => data_out <= "000";
            when "00011110000110" => data_out <= "000";
            when "00011110000111" => data_out <= "000";
            when "00011110001000" => data_out <= "000";
            when "00011110001001" => data_out <= "000";
            when "00011110001010" => data_out <= "000";
            when "00011110001011" => data_out <= "000";
            when "00011110001100" => data_out <= "000";
            when "00011110001101" => data_out <= "000";
            when "00011110001110" => data_out <= "000";
            when "00011110001111" => data_out <= "000";
            when "00011110010000" => data_out <= "000";
            when "00011110010001" => data_out <= "000";
            when "00011110010010" => data_out <= "000";
            when "00011110010011" => data_out <= "000";
            when "00011110010100" => data_out <= "000";
            when "00011110010101" => data_out <= "000";
            when "00011110010110" => data_out <= "000";
            when "00011110010111" => data_out <= "000";
            when "00011110011000" => data_out <= "000";
            when "00011110011001" => data_out <= "000";
            when "00011110011010" => data_out <= "000";
            when "00011110011011" => data_out <= "000";
            when "00011110011100" => data_out <= "000";
            when "00011110011101" => data_out <= "000";
            when "00011110011110" => data_out <= "000";
            when "00011110011111" => data_out <= "000";
            when "00011110100000" => data_out <= "000";
            when "00011110100001" => data_out <= "000";
            when "00011110100010" => data_out <= "000";
            when "00011110100011" => data_out <= "000";
            when "00011110100100" => data_out <= "000";
            when "00011110100101" => data_out <= "000";
            when "00011110100110" => data_out <= "000";
            when "00011110100111" => data_out <= "000";
            when "00011110101000" => data_out <= "000";
            when "00011110101001" => data_out <= "000";
            when "00011110101010" => data_out <= "000";
            when "00011110101011" => data_out <= "000";
            when "00011110101100" => data_out <= "000";
            when "00011110101101" => data_out <= "000";
            when "00011110101110" => data_out <= "000";
            when "00011110101111" => data_out <= "000";
            when "00011110110000" => data_out <= "000";
            when "00011110110001" => data_out <= "000";
            when "00011110110010" => data_out <= "000";
            when "00011110110011" => data_out <= "000";
            when "00011110110100" => data_out <= "000";
            when "00011110110101" => data_out <= "000";
            when "00011110110110" => data_out <= "000";
            when "00011110110111" => data_out <= "000";
            when "00011110111000" => data_out <= "000";
            when "00011110111001" => data_out <= "000";
            when "00011110111010" => data_out <= "000";
            when "00011110111011" => data_out <= "000";
            when "00011110111100" => data_out <= "000";
            when "00011110111101" => data_out <= "000";
            when "00011110111110" => data_out <= "000";
            when "00011110111111" => data_out <= "000";
            when "00011111000000" => data_out <= "000";
            when "00011111000001" => data_out <= "000";
            when "00011111000010" => data_out <= "000";
            when "00011111000011" => data_out <= "000";
            when "00011111000100" => data_out <= "000";
            when "00011111000101" => data_out <= "000";
            when "00011111000110" => data_out <= "000";
            when "00011111000111" => data_out <= "000";
            when "00011111001000" => data_out <= "000";
            when "00011111001001" => data_out <= "000";
            when "00011111001010" => data_out <= "000";
            when "00011111001011" => data_out <= "000";
            when "00011111001100" => data_out <= "000";
            when "00011111001101" => data_out <= "000";
            when "00011111001110" => data_out <= "000";
            when "00011111001111" => data_out <= "000";
            when "00011111010000" => data_out <= "000";
            when "00011111010001" => data_out <= "000";
            when "00011111010010" => data_out <= "000";
            when "00011111010011" => data_out <= "000";
            when "00011111010100" => data_out <= "000";
            when "00011111010101" => data_out <= "000";
            when "00011111010110" => data_out <= "000";
            when "00011111010111" => data_out <= "000";
            when "00011111011000" => data_out <= "000";
            when "00011111011001" => data_out <= "000";
            when "00011111011010" => data_out <= "000";
            when "00011111011011" => data_out <= "000";
            when "00011111011100" => data_out <= "000";
            when "00011111011101" => data_out <= "000";
            when "00011111011110" => data_out <= "000";
            when "00011111011111" => data_out <= "000";
            when "00011111100000" => data_out <= "000";
            when "00011111100001" => data_out <= "000";
            when "00011111100010" => data_out <= "000";
            when "00011111100011" => data_out <= "000";
            when "00011111100100" => data_out <= "000";
            when "00011111100101" => data_out <= "000";
            when "00011111100110" => data_out <= "000";
            when "00011111100111" => data_out <= "000";
            when "00011111101000" => data_out <= "000";
            when "00011111101001" => data_out <= "000";
            when "00011111101010" => data_out <= "000";
            when "00011111101011" => data_out <= "000";
            when "00011111101100" => data_out <= "000";
            when "00011111101101" => data_out <= "000";
            when "00011111101110" => data_out <= "000";
            when "00011111101111" => data_out <= "000";
            when "00011111110000" => data_out <= "000";
            when "00011111110001" => data_out <= "000";
            when "00011111110010" => data_out <= "000";
            when "00011111110011" => data_out <= "000";
            when "00011111110100" => data_out <= "000";
            when "00011111110101" => data_out <= "000";
            when "00011111110110" => data_out <= "000";
            when "00011111110111" => data_out <= "000";
            when "00011111111000" => data_out <= "000";
            when "00011111111001" => data_out <= "000";
            when "00011111111010" => data_out <= "000";
            when "00011111111011" => data_out <= "000";
            when "00011111111100" => data_out <= "000";
            when "00011111111101" => data_out <= "000";
            when "00011111111110" => data_out <= "000";
            when "00011111111111" => data_out <= "000";
            when others => data_out <= (others => '0'); -- Default case
        end case;
    end process;

end Behavioral;
